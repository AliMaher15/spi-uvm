package axi_item_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import axi_global_params_pkg::DATA_WIDTH;

    
    `include "axi_item_c.svh"
  
endpackage : axi_item_pkg