interface spi_slave_intf
                      (
                        input i_Clk,
                        input i_Rst_L
                      );

// Control/Data Signals
logic                         o_RX_DV;      // Data Valid pulse (1 clock cycle)                   
logic         [7:0]           o_RX_Byte;    // Byte received on MOSI
logic                         i_TX_DV;      // Data Valid pulse to register i_TX_Byte (by user)
logic         [7:0]           i_TX_Byte;    // Byte to serialize to MISO.             (by user)
// SPI Interface
logic                         i_SPI_Clk;    // slave clock generated by master (IDLE = 0 in mode 1)
logic                         o_SPI_MISO;   // master input, slave output serialized data (LSB first)
logic                         i_SPI_MOSI;   // master output, slave input serialized data (MSB first)
logic                         i_SPI_CS_n;   // active low, if this slave is selected to be active (controlled by higher logic)


//********* MACROS FUNCTIONS ***********//
`define spi_s_assert_clk(arg) \
  assert property (@(posedge CLK) disable iff (!RST) arg);

`define spi_s_assert_async_rst(arg) \
  assert property (@(negedge RST) 1'b1 |=> @(posedge CLK) arg);


Assert_SPI_Slave_MISO_is_tristate_when_CS_high :
  `spi_s_assert_clk(i_SPI_CS_n |-> o_SPI_MISO == 1'bz)
    
endinterface : spi_slave_intf