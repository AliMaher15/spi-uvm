package axi_global_params_pkg;

    parameter   CLK_PERIOD        = `def_axi_CLK_PERIOD;
    parameter   DATA_WIDTH        = `def_axi_DATA_WIDTH;
    
endpackage: axi_global_params_pkg