// Interface: spi_master_intf
//
interface spi_master_intf
                      (
                        input i_Clk,
                        input i_Rst_L
                      );

// TX (MOSI) Signals
logic    [7:0]    i_TX_Byte;        // Byte to transmit on MOSI
logic             i_TX_DV;          // Data Valid Pulse with i_TX_Byte
logic             o_TX_Ready;       // Transmit Ready for next byte

// RX (MISO) Signals
logic             o_RX_DV;          // Data Valid pulse (1 clock cycle)
logic    [7:0]    o_RX_Byte;        // Byte received on MISO

// SPI Interface
logic             i_SPI_MISO;       // master input, slave output serialized data (LSB first)
logic             o_SPI_MOSI;       // master output, slave input serialized data (MSB first)
logic             o_SPI_Clk;        // slave clock generated by master (at Mode "0"/"1" = 0)


//********* MACROS FUNCTIONS ***********//
`define spi_master_assert_clk(arg) \
  assert property (@(posedge CLK) disable iff (!RST) arg);

`define spi_master_assert_async_rst(arg) \
  assert property (@(negedge RST) 1'b1 |=> @(posedge CLK) arg);


Assert_spi_master_rst_control_signals :
  `spi_master_assert_async_rst(i_TX_Byte==0 && i_TX_DV==0 && o_TX_Ready==0 && o_RX_DV && o_RX_Byte)

Assert_spi_master_rst_interface_signals :
  `spi_master_assert_async_rst(i_SPI_MISO==0 && o_SPI_MOSI==0)
    
endinterface : spi_master_intf