interface rst_intf ();

    logic    res_n;    //output
    
endinterface : rst_intf