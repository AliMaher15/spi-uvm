// Interface: spi_master_intf
//
interface spi_master_intf
                      (
                        input i_Clk,
                        input i_Rst_L
                      );

// SPI Interface
logic             i_SPI_MISO;       // master input, slave output serialized data (LSB first)
logic             o_SPI_MOSI;       // master output, slave input serialized data (MSB first)
logic             o_SPI_Clk;        // slave clock generated by master (at Mode "0"/"1" = 0)


//********* MACROS FUNCTIONS ***********//
`define spi_master_assert_clk(arg) \
  assert property (@(posedge CLK) disable iff (!RST) arg);

`define spi_master_assert_async_rst(arg) \
  assert property (@(negedge RST) 1'b1 |=> @(posedge CLK) arg);


Assert_spi_master_rst_control_signals :
  `spi_master_assert_async_rst(i_TX_Byte==0 && i_TX_DV==0 && o_TX_Ready==0 && o_RX_DV && o_RX_Byte)

Assert_spi_master_rst_interface_signals :
  `spi_master_assert_async_rst(i_SPI_MISO==0 && o_SPI_MOSI==0)
    
endinterface : spi_master_intf