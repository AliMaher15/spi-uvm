package spi_seq_pkg ;
    
	import uvm_pkg::*;
	`include "uvm_macros.svh"

    import spi_item_pkg::*;
    import spi_tb_pkg::*;
    

    `include "spi_base_seq_c.svh"  
    `include "spi_general_seq_c.svh"
    `include "spi_gnrl_constr_seq_c.svh"

   

endpackage : spi_seq_pkg