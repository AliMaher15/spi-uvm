package spi_item_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    
    `include "spi_item_c.svh"
  
endpackage : spi_item_pkg