package spi_global_params_pkg;

    parameter   CLK_PERIOD        = `def_spi_CLK_PERIOD;
    
endpackage: spi_global_params_pkg