package axi_seq_pkg ;
    
	import uvm_pkg::*;
	`include "uvm_macros.svh"

    import axi_item_pkg::*;
    import axi_tb_pkg::*;
    

    `include "axi_base_seq_c.svh"  
           
    `include "axi_seq_c.svh"
    //`include "axi_master_seq_c.svh"
    //`include "axi_slave_seq_c.svh"
   

endpackage : axi_seq_pkg